
module SYS_TOP 
(
 input   wire                          RST_N,
 input   wire                          UART_CLK,
 input   wire                          REF_CLK,
 input   wire                          UART_RX_IN,
 output  wire                          UART_TX_O,
 output  wire                          parity_error,
 output  wire                          framing_error
);




///********************************************************///
//////////////////// Reset synchronizers /////////////////////
///********************************************************///




///********************************************************///
///////////////////// Data Synchronizers /////////////////////
///********************************************************///



///********************************************************///
///////////////////////// Async FIFO /////////////////////////
///********************************************************///



///********************************************************///
//////////////////////// Pulse Generator /////////////////////
///********************************************************///


///********************************************************///
//////////// Clock Divider for UART_TX Clock /////////////////
///********************************************************///



///********************************************************///
/////////////////////// Custom Mux Clock /////////////////////
///********************************************************///


///********************************************************///
//////////// Clock Divider for UART_RX Clock /////////////////
///********************************************************///



///********************************************************///
/////////////////////////// UART /////////////////////////////
///********************************************************///



///********************************************************///
//////////////////// System Controller ///////////////////////
///********************************************************///



///********************************************************///
/////////////////////// Register File ////////////////////////
///********************************************************///



///********************************************************///
//////////////////////////// ALU /////////////////////////////
///********************************************************///
 


///********************************************************///
///////////////////////// Clock Gating ///////////////////////
///********************************************************///




endmodule
 